module Top (
        input clk,
        nRst
    );
    
endmodule