module one_valid_16 (
    input  [15:0] in,
    output [ 3:0] out_en
);

wire [15:0] one_in;

assign one_in[0] = in[0];

genvar i;
generate 
	for (i=1; i<16; i=i+1)
	begin: sel_one
		assign one_in[i] = in[i] && ~|in[i-1:0];
	end
endgenerate

encoder_16_4 coder (.in(one_in), .out(out_en));

endmodule

module one_valid_32 (
    input  [31:0] in,
    output [ 4:0] out_en
);

wire [31:0] one_in;

assign one_in[0] = in[0];

genvar i;
generate 
	for (i=1; i<32; i=i+1)
	begin: sel_one
		assign one_in[i] = in[i] && ~|in[i-1:0];
	end
endgenerate

encoder_32_5 coder (.in(one_in), .out(out_en));

endmodule


module encoder_16_4(
    input  [15:0] in,
    output [ 3:0] out
);

wire [1:0] out_0, out_1, out_2, out_3;

encoder_4_2 one (.in(in[ 3: 0]), .out(out_0));
encoder_4_2 two (.in(in[ 7: 4]), .out(out_1));
encoder_4_2 thr (.in(in[11: 8]), .out(out_2));
encoder_4_2 fou (.in(in[15:12]), .out(out_3));

assign out = {4{|in[ 3: 0]}} & {2'd0, out_0} |
	     {4{|in[ 7: 4]}} & {2'd1, out_1} |		
	     {4{|in[11: 8]}} & {2'd2, out_2} |		
	     {4{|in[15:12]}} & {2'd3, out_3} ;		

endmodule


module encoder_32_5(
    input  [31:0] in,
    output [ 4:0] out
);

wire [3:0] out_0, out_1;

encoder_16_4 one (.in(in[15: 0]), .out(out_0));
encoder_16_4 two (.in(in[31:16]), .out(out_1));

assign out = {5{|in[15: 0]}} & {1'd0, out_0} |
	     {5{|in[31:16]}} & {1'd1, out_1} ;

endmodule

module decoder_2_4 (
    input wire [1:0] in,
    output reg [3:0] out
);
    always @ (*) begin
        case(in)
            2'b00:begin out = 4'b0001; end
            2'b01:begin out = 4'b0010; end
            2'b10:begin out = 4'b0100; end
            2'b11:begin out = 4'b1000; end
            default:begin
                out = 4'b0000;
            end
        endcase
    end
endmodule 



module decoder_3_8 (
    input wire [2:0] in,
    output reg [7:0] out
);
    always @ (*) begin
        case(in)
            3'b000:begin out = 8'b1; end
            3'b001:begin out = 8'b10; end
            3'b010:begin out = 8'b100; end
            3'b011:begin out = 8'b1000; end
            3'b100:begin out = 8'b10000; end
            3'b101:begin out = 8'b100000; end
            3'b110:begin out = 8'b1000000; end 
            3'b111:begin out = 8'b10000000; end
            default:begin
                out = 8'b0;
            end
        endcase
    end
endmodule 



module decoder_4_16(
    input wire [3:0] in,
    output reg [15:0] out
);
    always @ (*) begin
        case(in)
            4'd0:begin out = 16'b1; end
            4'd1:begin out = 16'b10; end
            4'd2:begin out = 16'b100; end
            4'd3:begin out = 16'b1000; end
            4'd4:begin out = 16'b10000; end
            4'd5:begin out = 16'b100000; end
            4'd6:begin out = 16'b1000000; end
            4'd7:begin out = 16'b10000000; end
            4'd8:begin out = 16'b100000000; end
            4'd9:begin out = 16'b1000000000; end
            4'd10:begin out = 16'b10000000000; end
            4'd11:begin out = 16'b100000000000; end
            4'd12:begin out = 16'b1000000000000; end
            4'd13:begin out = 16'b10000000000000; end
            4'd14:begin out = 16'b100000000000000; end
            4'd15:begin out = 16'b1000000000000000; end
            default:begin
                out = 16'b0;
            end
        endcase 
    end
endmodule



module decoder_5_32 (
    input wire [4:0] in,
    output reg [31:0] out
);
    always @ (*) begin
        case(in)
            5'd00:begin out=32'b00000000000000000000000000000001; end
            5'd01:begin out=32'b00000000000000000000000000000010; end
            5'd02:begin out=32'b00000000000000000000000000000100; end
            5'd03:begin out=32'b00000000000000000000000000001000; end
            5'd04:begin out=32'b00000000000000000000000000010000; end
            5'd05:begin out=32'b00000000000000000000000000100000; end
            5'd06:begin out=32'b00000000000000000000000001000000; end
            5'd07:begin out=32'b00000000000000000000000010000000; end
            5'd08:begin out=32'b00000000000000000000000100000000; end
            5'd09:begin out=32'b00000000000000000000001000000000; end
            5'd10:begin out=32'b00000000000000000000010000000000; end
            5'd11:begin out=32'b00000000000000000000100000000000; end
            5'd12:begin out=32'b00000000000000000001000000000000; end
            5'd13:begin out=32'b00000000000000000010000000000000; end
            5'd14:begin out=32'b00000000000000000100000000000000; end
            5'd15:begin out=32'b00000000000000001000000000000000; end
            5'd16:begin out=32'b00000000000000010000000000000000; end
            5'd17:begin out=32'b00000000000000100000000000000000; end
            5'd18:begin out=32'b00000000000001000000000000000000; end
            5'd19:begin out=32'b00000000000010000000000000000000; end
            5'd20:begin out=32'b00000000000100000000000000000000; end
            5'd21:begin out=32'b00000000001000000000000000000000; end
            5'd22:begin out=32'b00000000010000000000000000000000; end
            5'd23:begin out=32'b00000000100000000000000000000000; end
            5'd24:begin out=32'b00000001000000000000000000000000; end
            5'd25:begin out=32'b00000010000000000000000000000000; end
            5'd26:begin out=32'b00000100000000000000000000000000; end
            5'd27:begin out=32'b00001000000000000000000000000000; end
            5'd28:begin out=32'b00010000000000000000000000000000; end
            5'd29:begin out=32'b00100000000000000000000000000000; end
            5'd30:begin out=32'b01000000000000000000000000000000; end
            5'd31:begin out=32'b10000000000000000000000000000000; end
            default:begin
                out=32'b0;
            end
        endcase
    end
endmodule



module decoder_6_64 (
    input wire [5:0] in,
    output reg [63:0] out
);
    always @ (*) begin
        case(in)
            6'd00:begin out=64'b0000000000000000000000000000000000000000000000000000000000000001; end
            6'd01:begin out=64'b0000000000000000000000000000000000000000000000000000000000000010; end
            6'd02:begin out=64'b0000000000000000000000000000000000000000000000000000000000000100; end
            6'd03:begin out=64'b0000000000000000000000000000000000000000000000000000000000001000; end
            6'd04:begin out=64'b0000000000000000000000000000000000000000000000000000000000010000; end
            6'd05:begin out=64'b0000000000000000000000000000000000000000000000000000000000100000; end
            6'd06:begin out=64'b0000000000000000000000000000000000000000000000000000000001000000; end
            6'd07:begin out=64'b0000000000000000000000000000000000000000000000000000000010000000; end
            6'd08:begin out=64'b0000000000000000000000000000000000000000000000000000000100000000; end
            6'd09:begin out=64'b0000000000000000000000000000000000000000000000000000001000000000; end
            6'd10:begin out=64'b0000000000000000000000000000000000000000000000000000010000000000; end
            6'd11:begin out=64'b0000000000000000000000000000000000000000000000000000100000000000; end
            6'd12:begin out=64'b0000000000000000000000000000000000000000000000000001000000000000; end
            6'd13:begin out=64'b0000000000000000000000000000000000000000000000000010000000000000; end
            6'd14:begin out=64'b0000000000000000000000000000000000000000000000000100000000000000; end
            6'd15:begin out=64'b0000000000000000000000000000000000000000000000001000000000000000; end
            6'd16:begin out=64'b0000000000000000000000000000000000000000000000010000000000000000; end
            6'd17:begin out=64'b0000000000000000000000000000000000000000000000100000000000000000; end
            6'd18:begin out=64'b0000000000000000000000000000000000000000000001000000000000000000; end
            6'd19:begin out=64'b0000000000000000000000000000000000000000000010000000000000000000; end
            6'd20:begin out=64'b0000000000000000000000000000000000000000000100000000000000000000; end
            6'd21:begin out=64'b0000000000000000000000000000000000000000001000000000000000000000; end
            6'd22:begin out=64'b0000000000000000000000000000000000000000010000000000000000000000; end
            6'd23:begin out=64'b0000000000000000000000000000000000000000100000000000000000000000; end
            6'd24:begin out=64'b0000000000000000000000000000000000000001000000000000000000000000; end
            6'd25:begin out=64'b0000000000000000000000000000000000000010000000000000000000000000; end
            6'd26:begin out=64'b0000000000000000000000000000000000000100000000000000000000000000; end
            6'd27:begin out=64'b0000000000000000000000000000000000001000000000000000000000000000; end
            6'd28:begin out=64'b0000000000000000000000000000000000010000000000000000000000000000; end
            6'd29:begin out=64'b0000000000000000000000000000000000100000000000000000000000000000; end
            6'd30:begin out=64'b0000000000000000000000000000000001000000000000000000000000000000; end
            6'd31:begin out=64'b0000000000000000000000000000000010000000000000000000000000000000; end
            6'd32:begin out=64'b0000000000000000000000000000000100000000000000000000000000000000; end
            6'd33:begin out=64'b0000000000000000000000000000001000000000000000000000000000000000; end
            6'd34:begin out=64'b0000000000000000000000000000010000000000000000000000000000000000; end
            6'd35:begin out=64'b0000000000000000000000000000100000000000000000000000000000000000; end
            6'd36:begin out=64'b0000000000000000000000000001000000000000000000000000000000000000; end
            6'd37:begin out=64'b0000000000000000000000000010000000000000000000000000000000000000; end
            6'd38:begin out=64'b0000000000000000000000000100000000000000000000000000000000000000; end
            6'd39:begin out=64'b0000000000000000000000001000000000000000000000000000000000000000; end
            6'd40:begin out=64'b0000000000000000000000010000000000000000000000000000000000000000; end
            6'd41:begin out=64'b0000000000000000000000100000000000000000000000000000000000000000; end
            6'd42:begin out=64'b0000000000000000000001000000000000000000000000000000000000000000; end
            6'd43:begin out=64'b0000000000000000000010000000000000000000000000000000000000000000; end
            6'd44:begin out=64'b0000000000000000000100000000000000000000000000000000000000000000; end
            6'd45:begin out=64'b0000000000000000001000000000000000000000000000000000000000000000; end
            6'd46:begin out=64'b0000000000000000010000000000000000000000000000000000000000000000; end
            6'd47:begin out=64'b0000000000000000100000000000000000000000000000000000000000000000; end
            6'd48:begin out=64'b0000000000000001000000000000000000000000000000000000000000000000; end
            6'd49:begin out=64'b0000000000000010000000000000000000000000000000000000000000000000; end
            6'd50:begin out=64'b0000000000000100000000000000000000000000000000000000000000000000; end
            6'd51:begin out=64'b0000000000001000000000000000000000000000000000000000000000000000; end
            6'd52:begin out=64'b0000000000010000000000000000000000000000000000000000000000000000; end
            6'd53:begin out=64'b0000000000100000000000000000000000000000000000000000000000000000; end
            6'd54:begin out=64'b0000000001000000000000000000000000000000000000000000000000000000; end
            6'd55:begin out=64'b0000000010000000000000000000000000000000000000000000000000000000; end
            6'd56:begin out=64'b0000000100000000000000000000000000000000000000000000000000000000; end
            6'd57:begin out=64'b0000001000000000000000000000000000000000000000000000000000000000; end
            6'd58:begin out=64'b0000010000000000000000000000000000000000000000000000000000000000; end
            6'd59:begin out=64'b0000100000000000000000000000000000000000000000000000000000000000; end
            6'd60:begin out=64'b0001000000000000000000000000000000000000000000000000000000000000; end
            6'd61:begin out=64'b0010000000000000000000000000000000000000000000000000000000000000; end
            6'd62:begin out=64'b0100000000000000000000000000000000000000000000000000000000000000; end
            6'd63:begin out=64'b1000000000000000000000000000000000000000000000000000000000000000; end   
            default:begin
                out=64'b0;
            end
        endcase
    end

endmodule 