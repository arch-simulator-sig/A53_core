module decoder_5_32 (
    input wire [4:0] in,
    output reg [31:0] out
);
    always @ (*) begin
        case(in)
            5'd00:begin out=32'b00000000000000000000000000000001; end
            5'd01:begin out=32'b00000000000000000000000000000010; end
            5'd02:begin out=32'b00000000000000000000000000000100; end
            5'd03:begin out=32'b00000000000000000000000000001000; end
            5'd04:begin out=32'b00000000000000000000000000010000; end
            5'd05:begin out=32'b00000000000000000000000000100000; end
            5'd06:begin out=32'b00000000000000000000000001000000; end
            5'd07:begin out=32'b00000000000000000000000010000000; end
            5'd08:begin out=32'b00000000000000000000000100000000; end
            5'd09:begin out=32'b00000000000000000000001000000000; end
            5'd10:begin out=32'b00000000000000000000010000000000; end
            5'd11:begin out=32'b00000000000000000000100000000000; end
            5'd12:begin out=32'b00000000000000000001000000000000; end
            5'd13:begin out=32'b00000000000000000010000000000000; end
            5'd14:begin out=32'b00000000000000000100000000000000; end
            5'd15:begin out=32'b00000000000000001000000000000000; end
            5'd16:begin out=32'b00000000000000010000000000000000; end
            5'd17:begin out=32'b00000000000000100000000000000000; end
            5'd18:begin out=32'b00000000000001000000000000000000; end
            5'd19:begin out=32'b00000000000010000000000000000000; end
            5'd20:begin out=32'b00000000000100000000000000000000; end
            5'd21:begin out=32'b00000000001000000000000000000000; end
            5'd22:begin out=32'b00000000010000000000000000000000; end
            5'd23:begin out=32'b00000000100000000000000000000000; end
            5'd24:begin out=32'b00000001000000000000000000000000; end
            5'd25:begin out=32'b00000010000000000000000000000000; end
            5'd26:begin out=32'b00000100000000000000000000000000; end
            5'd27:begin out=32'b00001000000000000000000000000000; end
            5'd28:begin out=32'b00010000000000000000000000000000; end
            5'd29:begin out=32'b00100000000000000000000000000000; end
            5'd30:begin out=32'b01000000000000000000000000000000; end
            5'd31:begin out=32'b10000000000000000000000000000000; end
            default:begin
                out=32'b0;
            end
        endcase
    end
endmodule